magic
tech sky130B
magscale 1 2
timestamp 1686588514
<< pwell >>
rect -1457 -1319 1457 1319
<< nmoslvt >>
rect -1261 109 -1061 1109
rect -1003 109 -803 1109
rect -745 109 -545 1109
rect -487 109 -287 1109
rect -229 109 -29 1109
rect 29 109 229 1109
rect 287 109 487 1109
rect 545 109 745 1109
rect 803 109 1003 1109
rect 1061 109 1261 1109
rect -1261 -1109 -1061 -109
rect -1003 -1109 -803 -109
rect -745 -1109 -545 -109
rect -487 -1109 -287 -109
rect -229 -1109 -29 -109
rect 29 -1109 229 -109
rect 287 -1109 487 -109
rect 545 -1109 745 -109
rect 803 -1109 1003 -109
rect 1061 -1109 1261 -109
<< ndiff >>
rect -1319 1097 -1261 1109
rect -1319 121 -1307 1097
rect -1273 121 -1261 1097
rect -1319 109 -1261 121
rect -1061 1097 -1003 1109
rect -1061 121 -1049 1097
rect -1015 121 -1003 1097
rect -1061 109 -1003 121
rect -803 1097 -745 1109
rect -803 121 -791 1097
rect -757 121 -745 1097
rect -803 109 -745 121
rect -545 1097 -487 1109
rect -545 121 -533 1097
rect -499 121 -487 1097
rect -545 109 -487 121
rect -287 1097 -229 1109
rect -287 121 -275 1097
rect -241 121 -229 1097
rect -287 109 -229 121
rect -29 1097 29 1109
rect -29 121 -17 1097
rect 17 121 29 1097
rect -29 109 29 121
rect 229 1097 287 1109
rect 229 121 241 1097
rect 275 121 287 1097
rect 229 109 287 121
rect 487 1097 545 1109
rect 487 121 499 1097
rect 533 121 545 1097
rect 487 109 545 121
rect 745 1097 803 1109
rect 745 121 757 1097
rect 791 121 803 1097
rect 745 109 803 121
rect 1003 1097 1061 1109
rect 1003 121 1015 1097
rect 1049 121 1061 1097
rect 1003 109 1061 121
rect 1261 1097 1319 1109
rect 1261 121 1273 1097
rect 1307 121 1319 1097
rect 1261 109 1319 121
rect -1319 -121 -1261 -109
rect -1319 -1097 -1307 -121
rect -1273 -1097 -1261 -121
rect -1319 -1109 -1261 -1097
rect -1061 -121 -1003 -109
rect -1061 -1097 -1049 -121
rect -1015 -1097 -1003 -121
rect -1061 -1109 -1003 -1097
rect -803 -121 -745 -109
rect -803 -1097 -791 -121
rect -757 -1097 -745 -121
rect -803 -1109 -745 -1097
rect -545 -121 -487 -109
rect -545 -1097 -533 -121
rect -499 -1097 -487 -121
rect -545 -1109 -487 -1097
rect -287 -121 -229 -109
rect -287 -1097 -275 -121
rect -241 -1097 -229 -121
rect -287 -1109 -229 -1097
rect -29 -121 29 -109
rect -29 -1097 -17 -121
rect 17 -1097 29 -121
rect -29 -1109 29 -1097
rect 229 -121 287 -109
rect 229 -1097 241 -121
rect 275 -1097 287 -121
rect 229 -1109 287 -1097
rect 487 -121 545 -109
rect 487 -1097 499 -121
rect 533 -1097 545 -121
rect 487 -1109 545 -1097
rect 745 -121 803 -109
rect 745 -1097 757 -121
rect 791 -1097 803 -121
rect 745 -1109 803 -1097
rect 1003 -121 1061 -109
rect 1003 -1097 1015 -121
rect 1049 -1097 1061 -121
rect 1003 -1109 1061 -1097
rect 1261 -121 1319 -109
rect 1261 -1097 1273 -121
rect 1307 -1097 1319 -121
rect 1261 -1109 1319 -1097
<< ndiffc >>
rect -1307 121 -1273 1097
rect -1049 121 -1015 1097
rect -791 121 -757 1097
rect -533 121 -499 1097
rect -275 121 -241 1097
rect -17 121 17 1097
rect 241 121 275 1097
rect 499 121 533 1097
rect 757 121 791 1097
rect 1015 121 1049 1097
rect 1273 121 1307 1097
rect -1307 -1097 -1273 -121
rect -1049 -1097 -1015 -121
rect -791 -1097 -757 -121
rect -533 -1097 -499 -121
rect -275 -1097 -241 -121
rect -17 -1097 17 -121
rect 241 -1097 275 -121
rect 499 -1097 533 -121
rect 757 -1097 791 -121
rect 1015 -1097 1049 -121
rect 1273 -1097 1307 -121
<< psubdiff >>
rect -1421 1249 -1325 1283
rect 1325 1249 1421 1283
rect -1421 1187 -1387 1249
rect 1387 1187 1421 1249
rect -1421 -1249 -1387 -1187
rect 1387 -1249 1421 -1187
rect -1421 -1283 -1325 -1249
rect 1325 -1283 1421 -1249
<< psubdiffcont >>
rect -1325 1249 1325 1283
rect -1421 -1187 -1387 1187
rect 1387 -1187 1421 1187
rect -1325 -1283 1325 -1249
<< poly >>
rect -1227 1181 -1095 1197
rect -1227 1164 -1211 1181
rect -1261 1147 -1211 1164
rect -1111 1164 -1095 1181
rect -969 1181 -837 1197
rect -969 1164 -953 1181
rect -1111 1147 -1061 1164
rect -1261 1109 -1061 1147
rect -1003 1147 -953 1164
rect -853 1164 -837 1181
rect -711 1181 -579 1197
rect -711 1164 -695 1181
rect -853 1147 -803 1164
rect -1003 1109 -803 1147
rect -745 1147 -695 1164
rect -595 1164 -579 1181
rect -453 1181 -321 1197
rect -453 1164 -437 1181
rect -595 1147 -545 1164
rect -745 1109 -545 1147
rect -487 1147 -437 1164
rect -337 1164 -321 1181
rect -195 1181 -63 1197
rect -195 1164 -179 1181
rect -337 1147 -287 1164
rect -487 1109 -287 1147
rect -229 1147 -179 1164
rect -79 1164 -63 1181
rect 63 1181 195 1197
rect 63 1164 79 1181
rect -79 1147 -29 1164
rect -229 1109 -29 1147
rect 29 1147 79 1164
rect 179 1164 195 1181
rect 321 1181 453 1197
rect 321 1164 337 1181
rect 179 1147 229 1164
rect 29 1109 229 1147
rect 287 1147 337 1164
rect 437 1164 453 1181
rect 579 1181 711 1197
rect 579 1164 595 1181
rect 437 1147 487 1164
rect 287 1109 487 1147
rect 545 1147 595 1164
rect 695 1164 711 1181
rect 837 1181 969 1197
rect 837 1164 853 1181
rect 695 1147 745 1164
rect 545 1109 745 1147
rect 803 1147 853 1164
rect 953 1164 969 1181
rect 1095 1181 1227 1197
rect 1095 1164 1111 1181
rect 953 1147 1003 1164
rect 803 1109 1003 1147
rect 1061 1147 1111 1164
rect 1211 1164 1227 1181
rect 1211 1147 1261 1164
rect 1061 1109 1261 1147
rect -1261 71 -1061 109
rect -1261 54 -1211 71
rect -1227 37 -1211 54
rect -1111 54 -1061 71
rect -1003 71 -803 109
rect -1003 54 -953 71
rect -1111 37 -1095 54
rect -1227 21 -1095 37
rect -969 37 -953 54
rect -853 54 -803 71
rect -745 71 -545 109
rect -745 54 -695 71
rect -853 37 -837 54
rect -969 21 -837 37
rect -711 37 -695 54
rect -595 54 -545 71
rect -487 71 -287 109
rect -487 54 -437 71
rect -595 37 -579 54
rect -711 21 -579 37
rect -453 37 -437 54
rect -337 54 -287 71
rect -229 71 -29 109
rect -229 54 -179 71
rect -337 37 -321 54
rect -453 21 -321 37
rect -195 37 -179 54
rect -79 54 -29 71
rect 29 71 229 109
rect 29 54 79 71
rect -79 37 -63 54
rect -195 21 -63 37
rect 63 37 79 54
rect 179 54 229 71
rect 287 71 487 109
rect 287 54 337 71
rect 179 37 195 54
rect 63 21 195 37
rect 321 37 337 54
rect 437 54 487 71
rect 545 71 745 109
rect 545 54 595 71
rect 437 37 453 54
rect 321 21 453 37
rect 579 37 595 54
rect 695 54 745 71
rect 803 71 1003 109
rect 803 54 853 71
rect 695 37 711 54
rect 579 21 711 37
rect 837 37 853 54
rect 953 54 1003 71
rect 1061 71 1261 109
rect 1061 54 1111 71
rect 953 37 969 54
rect 837 21 969 37
rect 1095 37 1111 54
rect 1211 54 1261 71
rect 1211 37 1227 54
rect 1095 21 1227 37
rect -1227 -37 -1095 -21
rect -1227 -54 -1211 -37
rect -1261 -71 -1211 -54
rect -1111 -54 -1095 -37
rect -969 -37 -837 -21
rect -969 -54 -953 -37
rect -1111 -71 -1061 -54
rect -1261 -109 -1061 -71
rect -1003 -71 -953 -54
rect -853 -54 -837 -37
rect -711 -37 -579 -21
rect -711 -54 -695 -37
rect -853 -71 -803 -54
rect -1003 -109 -803 -71
rect -745 -71 -695 -54
rect -595 -54 -579 -37
rect -453 -37 -321 -21
rect -453 -54 -437 -37
rect -595 -71 -545 -54
rect -745 -109 -545 -71
rect -487 -71 -437 -54
rect -337 -54 -321 -37
rect -195 -37 -63 -21
rect -195 -54 -179 -37
rect -337 -71 -287 -54
rect -487 -109 -287 -71
rect -229 -71 -179 -54
rect -79 -54 -63 -37
rect 63 -37 195 -21
rect 63 -54 79 -37
rect -79 -71 -29 -54
rect -229 -109 -29 -71
rect 29 -71 79 -54
rect 179 -54 195 -37
rect 321 -37 453 -21
rect 321 -54 337 -37
rect 179 -71 229 -54
rect 29 -109 229 -71
rect 287 -71 337 -54
rect 437 -54 453 -37
rect 579 -37 711 -21
rect 579 -54 595 -37
rect 437 -71 487 -54
rect 287 -109 487 -71
rect 545 -71 595 -54
rect 695 -54 711 -37
rect 837 -37 969 -21
rect 837 -54 853 -37
rect 695 -71 745 -54
rect 545 -109 745 -71
rect 803 -71 853 -54
rect 953 -54 969 -37
rect 1095 -37 1227 -21
rect 1095 -54 1111 -37
rect 953 -71 1003 -54
rect 803 -109 1003 -71
rect 1061 -71 1111 -54
rect 1211 -54 1227 -37
rect 1211 -71 1261 -54
rect 1061 -109 1261 -71
rect -1261 -1147 -1061 -1109
rect -1261 -1164 -1211 -1147
rect -1227 -1181 -1211 -1164
rect -1111 -1164 -1061 -1147
rect -1003 -1147 -803 -1109
rect -1003 -1164 -953 -1147
rect -1111 -1181 -1095 -1164
rect -1227 -1197 -1095 -1181
rect -969 -1181 -953 -1164
rect -853 -1164 -803 -1147
rect -745 -1147 -545 -1109
rect -745 -1164 -695 -1147
rect -853 -1181 -837 -1164
rect -969 -1197 -837 -1181
rect -711 -1181 -695 -1164
rect -595 -1164 -545 -1147
rect -487 -1147 -287 -1109
rect -487 -1164 -437 -1147
rect -595 -1181 -579 -1164
rect -711 -1197 -579 -1181
rect -453 -1181 -437 -1164
rect -337 -1164 -287 -1147
rect -229 -1147 -29 -1109
rect -229 -1164 -179 -1147
rect -337 -1181 -321 -1164
rect -453 -1197 -321 -1181
rect -195 -1181 -179 -1164
rect -79 -1164 -29 -1147
rect 29 -1147 229 -1109
rect 29 -1164 79 -1147
rect -79 -1181 -63 -1164
rect -195 -1197 -63 -1181
rect 63 -1181 79 -1164
rect 179 -1164 229 -1147
rect 287 -1147 487 -1109
rect 287 -1164 337 -1147
rect 179 -1181 195 -1164
rect 63 -1197 195 -1181
rect 321 -1181 337 -1164
rect 437 -1164 487 -1147
rect 545 -1147 745 -1109
rect 545 -1164 595 -1147
rect 437 -1181 453 -1164
rect 321 -1197 453 -1181
rect 579 -1181 595 -1164
rect 695 -1164 745 -1147
rect 803 -1147 1003 -1109
rect 803 -1164 853 -1147
rect 695 -1181 711 -1164
rect 579 -1197 711 -1181
rect 837 -1181 853 -1164
rect 953 -1164 1003 -1147
rect 1061 -1147 1261 -1109
rect 1061 -1164 1111 -1147
rect 953 -1181 969 -1164
rect 837 -1197 969 -1181
rect 1095 -1181 1111 -1164
rect 1211 -1164 1261 -1147
rect 1211 -1181 1227 -1164
rect 1095 -1197 1227 -1181
<< polycont >>
rect -1211 1147 -1111 1181
rect -953 1147 -853 1181
rect -695 1147 -595 1181
rect -437 1147 -337 1181
rect -179 1147 -79 1181
rect 79 1147 179 1181
rect 337 1147 437 1181
rect 595 1147 695 1181
rect 853 1147 953 1181
rect 1111 1147 1211 1181
rect -1211 37 -1111 71
rect -953 37 -853 71
rect -695 37 -595 71
rect -437 37 -337 71
rect -179 37 -79 71
rect 79 37 179 71
rect 337 37 437 71
rect 595 37 695 71
rect 853 37 953 71
rect 1111 37 1211 71
rect -1211 -71 -1111 -37
rect -953 -71 -853 -37
rect -695 -71 -595 -37
rect -437 -71 -337 -37
rect -179 -71 -79 -37
rect 79 -71 179 -37
rect 337 -71 437 -37
rect 595 -71 695 -37
rect 853 -71 953 -37
rect 1111 -71 1211 -37
rect -1211 -1181 -1111 -1147
rect -953 -1181 -853 -1147
rect -695 -1181 -595 -1147
rect -437 -1181 -337 -1147
rect -179 -1181 -79 -1147
rect 79 -1181 179 -1147
rect 337 -1181 437 -1147
rect 595 -1181 695 -1147
rect 853 -1181 953 -1147
rect 1111 -1181 1211 -1147
<< locali >>
rect -1421 1249 -1325 1283
rect 1325 1249 1421 1283
rect -1421 1187 -1387 1249
rect 1387 1187 1421 1249
rect -1227 1147 -1211 1181
rect -1111 1147 -1095 1181
rect -969 1147 -953 1181
rect -853 1147 -837 1181
rect -711 1147 -695 1181
rect -595 1147 -579 1181
rect -453 1147 -437 1181
rect -337 1147 -321 1181
rect -195 1147 -179 1181
rect -79 1147 -63 1181
rect 63 1147 79 1181
rect 179 1147 195 1181
rect 321 1147 337 1181
rect 437 1147 453 1181
rect 579 1147 595 1181
rect 695 1147 711 1181
rect 837 1147 853 1181
rect 953 1147 969 1181
rect 1095 1147 1111 1181
rect 1211 1147 1227 1181
rect -1307 1097 -1273 1113
rect -1307 105 -1273 121
rect -1049 1097 -1015 1113
rect -1049 105 -1015 121
rect -791 1097 -757 1113
rect -791 105 -757 121
rect -533 1097 -499 1113
rect -533 105 -499 121
rect -275 1097 -241 1113
rect -275 105 -241 121
rect -17 1097 17 1113
rect -17 105 17 121
rect 241 1097 275 1113
rect 241 105 275 121
rect 499 1097 533 1113
rect 499 105 533 121
rect 757 1097 791 1113
rect 757 105 791 121
rect 1015 1097 1049 1113
rect 1015 105 1049 121
rect 1273 1097 1307 1113
rect 1273 105 1307 121
rect -1227 37 -1211 71
rect -1111 37 -1095 71
rect -969 37 -953 71
rect -853 37 -837 71
rect -711 37 -695 71
rect -595 37 -579 71
rect -453 37 -437 71
rect -337 37 -321 71
rect -195 37 -179 71
rect -79 37 -63 71
rect 63 37 79 71
rect 179 37 195 71
rect 321 37 337 71
rect 437 37 453 71
rect 579 37 595 71
rect 695 37 711 71
rect 837 37 853 71
rect 953 37 969 71
rect 1095 37 1111 71
rect 1211 37 1227 71
rect -1227 -71 -1211 -37
rect -1111 -71 -1095 -37
rect -969 -71 -953 -37
rect -853 -71 -837 -37
rect -711 -71 -695 -37
rect -595 -71 -579 -37
rect -453 -71 -437 -37
rect -337 -71 -321 -37
rect -195 -71 -179 -37
rect -79 -71 -63 -37
rect 63 -71 79 -37
rect 179 -71 195 -37
rect 321 -71 337 -37
rect 437 -71 453 -37
rect 579 -71 595 -37
rect 695 -71 711 -37
rect 837 -71 853 -37
rect 953 -71 969 -37
rect 1095 -71 1111 -37
rect 1211 -71 1227 -37
rect -1307 -121 -1273 -105
rect -1307 -1113 -1273 -1097
rect -1049 -121 -1015 -105
rect -1049 -1113 -1015 -1097
rect -791 -121 -757 -105
rect -791 -1113 -757 -1097
rect -533 -121 -499 -105
rect -533 -1113 -499 -1097
rect -275 -121 -241 -105
rect -275 -1113 -241 -1097
rect -17 -121 17 -105
rect -17 -1113 17 -1097
rect 241 -121 275 -105
rect 241 -1113 275 -1097
rect 499 -121 533 -105
rect 499 -1113 533 -1097
rect 757 -121 791 -105
rect 757 -1113 791 -1097
rect 1015 -121 1049 -105
rect 1015 -1113 1049 -1097
rect 1273 -121 1307 -105
rect 1273 -1113 1307 -1097
rect -1227 -1181 -1211 -1147
rect -1111 -1181 -1095 -1147
rect -969 -1181 -953 -1147
rect -853 -1181 -837 -1147
rect -711 -1181 -695 -1147
rect -595 -1181 -579 -1147
rect -453 -1181 -437 -1147
rect -337 -1181 -321 -1147
rect -195 -1181 -179 -1147
rect -79 -1181 -63 -1147
rect 63 -1181 79 -1147
rect 179 -1181 195 -1147
rect 321 -1181 337 -1147
rect 437 -1181 453 -1147
rect 579 -1181 595 -1147
rect 695 -1181 711 -1147
rect 837 -1181 853 -1147
rect 953 -1181 969 -1147
rect 1095 -1181 1111 -1147
rect 1211 -1181 1227 -1147
rect -1421 -1249 -1387 -1187
rect 1387 -1249 1421 -1187
rect -1421 -1283 -1325 -1249
rect 1325 -1283 1421 -1249
<< viali >>
rect -1211 1147 -1111 1181
rect -953 1147 -853 1181
rect -695 1147 -595 1181
rect -437 1147 -337 1181
rect -179 1147 -79 1181
rect 79 1147 179 1181
rect 337 1147 437 1181
rect 595 1147 695 1181
rect 853 1147 953 1181
rect 1111 1147 1211 1181
rect -1307 121 -1273 1097
rect -1049 121 -1015 1097
rect -791 121 -757 1097
rect -533 121 -499 1097
rect -275 121 -241 1097
rect -17 121 17 1097
rect 241 121 275 1097
rect 499 121 533 1097
rect 757 121 791 1097
rect 1015 121 1049 1097
rect 1273 121 1307 1097
rect -1211 37 -1111 71
rect -953 37 -853 71
rect -695 37 -595 71
rect -437 37 -337 71
rect -179 37 -79 71
rect 79 37 179 71
rect 337 37 437 71
rect 595 37 695 71
rect 853 37 953 71
rect 1111 37 1211 71
rect -1211 -71 -1111 -37
rect -953 -71 -853 -37
rect -695 -71 -595 -37
rect -437 -71 -337 -37
rect -179 -71 -79 -37
rect 79 -71 179 -37
rect 337 -71 437 -37
rect 595 -71 695 -37
rect 853 -71 953 -37
rect 1111 -71 1211 -37
rect -1307 -1097 -1273 -121
rect -1049 -1097 -1015 -121
rect -791 -1097 -757 -121
rect -533 -1097 -499 -121
rect -275 -1097 -241 -121
rect -17 -1097 17 -121
rect 241 -1097 275 -121
rect 499 -1097 533 -121
rect 757 -1097 791 -121
rect 1015 -1097 1049 -121
rect 1273 -1097 1307 -121
rect -1211 -1181 -1111 -1147
rect -953 -1181 -853 -1147
rect -695 -1181 -595 -1147
rect -437 -1181 -337 -1147
rect -179 -1181 -79 -1147
rect 79 -1181 179 -1147
rect 337 -1181 437 -1147
rect 595 -1181 695 -1147
rect 853 -1181 953 -1147
rect 1111 -1181 1211 -1147
<< metal1 >>
rect -1223 1181 -1099 1187
rect -1223 1147 -1211 1181
rect -1111 1147 -1099 1181
rect -1223 1141 -1099 1147
rect -965 1181 -841 1187
rect -965 1147 -953 1181
rect -853 1147 -841 1181
rect -965 1141 -841 1147
rect -707 1181 -583 1187
rect -707 1147 -695 1181
rect -595 1147 -583 1181
rect -707 1141 -583 1147
rect -449 1181 -325 1187
rect -449 1147 -437 1181
rect -337 1147 -325 1181
rect -449 1141 -325 1147
rect -191 1181 -67 1187
rect -191 1147 -179 1181
rect -79 1147 -67 1181
rect -191 1141 -67 1147
rect 67 1181 191 1187
rect 67 1147 79 1181
rect 179 1147 191 1181
rect 67 1141 191 1147
rect 325 1181 449 1187
rect 325 1147 337 1181
rect 437 1147 449 1181
rect 325 1141 449 1147
rect 583 1181 707 1187
rect 583 1147 595 1181
rect 695 1147 707 1181
rect 583 1141 707 1147
rect 841 1181 965 1187
rect 841 1147 853 1181
rect 953 1147 965 1181
rect 841 1141 965 1147
rect 1099 1181 1223 1187
rect 1099 1147 1111 1181
rect 1211 1147 1223 1181
rect 1099 1141 1223 1147
rect -1313 1097 -1267 1109
rect -1313 121 -1307 1097
rect -1273 121 -1267 1097
rect -1313 109 -1267 121
rect -1055 1097 -1009 1109
rect -1055 121 -1049 1097
rect -1015 121 -1009 1097
rect -1055 109 -1009 121
rect -797 1097 -751 1109
rect -797 121 -791 1097
rect -757 121 -751 1097
rect -797 109 -751 121
rect -539 1097 -493 1109
rect -539 121 -533 1097
rect -499 121 -493 1097
rect -539 109 -493 121
rect -281 1097 -235 1109
rect -281 121 -275 1097
rect -241 121 -235 1097
rect -281 109 -235 121
rect -23 1097 23 1109
rect -23 121 -17 1097
rect 17 121 23 1097
rect -23 109 23 121
rect 235 1097 281 1109
rect 235 121 241 1097
rect 275 121 281 1097
rect 235 109 281 121
rect 493 1097 539 1109
rect 493 121 499 1097
rect 533 121 539 1097
rect 493 109 539 121
rect 751 1097 797 1109
rect 751 121 757 1097
rect 791 121 797 1097
rect 751 109 797 121
rect 1009 1097 1055 1109
rect 1009 121 1015 1097
rect 1049 121 1055 1097
rect 1009 109 1055 121
rect 1267 1097 1313 1109
rect 1267 121 1273 1097
rect 1307 121 1313 1097
rect 1267 109 1313 121
rect -1223 71 -1099 77
rect -1223 37 -1211 71
rect -1111 37 -1099 71
rect -1223 31 -1099 37
rect -965 71 -841 77
rect -965 37 -953 71
rect -853 37 -841 71
rect -965 31 -841 37
rect -707 71 -583 77
rect -707 37 -695 71
rect -595 37 -583 71
rect -707 31 -583 37
rect -449 71 -325 77
rect -449 37 -437 71
rect -337 37 -325 71
rect -449 31 -325 37
rect -191 71 -67 77
rect -191 37 -179 71
rect -79 37 -67 71
rect -191 31 -67 37
rect 67 71 191 77
rect 67 37 79 71
rect 179 37 191 71
rect 67 31 191 37
rect 325 71 449 77
rect 325 37 337 71
rect 437 37 449 71
rect 325 31 449 37
rect 583 71 707 77
rect 583 37 595 71
rect 695 37 707 71
rect 583 31 707 37
rect 841 71 965 77
rect 841 37 853 71
rect 953 37 965 71
rect 841 31 965 37
rect 1099 71 1223 77
rect 1099 37 1111 71
rect 1211 37 1223 71
rect 1099 31 1223 37
rect -1223 -37 -1099 -31
rect -1223 -71 -1211 -37
rect -1111 -71 -1099 -37
rect -1223 -77 -1099 -71
rect -965 -37 -841 -31
rect -965 -71 -953 -37
rect -853 -71 -841 -37
rect -965 -77 -841 -71
rect -707 -37 -583 -31
rect -707 -71 -695 -37
rect -595 -71 -583 -37
rect -707 -77 -583 -71
rect -449 -37 -325 -31
rect -449 -71 -437 -37
rect -337 -71 -325 -37
rect -449 -77 -325 -71
rect -191 -37 -67 -31
rect -191 -71 -179 -37
rect -79 -71 -67 -37
rect -191 -77 -67 -71
rect 67 -37 191 -31
rect 67 -71 79 -37
rect 179 -71 191 -37
rect 67 -77 191 -71
rect 325 -37 449 -31
rect 325 -71 337 -37
rect 437 -71 449 -37
rect 325 -77 449 -71
rect 583 -37 707 -31
rect 583 -71 595 -37
rect 695 -71 707 -37
rect 583 -77 707 -71
rect 841 -37 965 -31
rect 841 -71 853 -37
rect 953 -71 965 -37
rect 841 -77 965 -71
rect 1099 -37 1223 -31
rect 1099 -71 1111 -37
rect 1211 -71 1223 -37
rect 1099 -77 1223 -71
rect -1313 -121 -1267 -109
rect -1313 -1097 -1307 -121
rect -1273 -1097 -1267 -121
rect -1313 -1109 -1267 -1097
rect -1055 -121 -1009 -109
rect -1055 -1097 -1049 -121
rect -1015 -1097 -1009 -121
rect -1055 -1109 -1009 -1097
rect -797 -121 -751 -109
rect -797 -1097 -791 -121
rect -757 -1097 -751 -121
rect -797 -1109 -751 -1097
rect -539 -121 -493 -109
rect -539 -1097 -533 -121
rect -499 -1097 -493 -121
rect -539 -1109 -493 -1097
rect -281 -121 -235 -109
rect -281 -1097 -275 -121
rect -241 -1097 -235 -121
rect -281 -1109 -235 -1097
rect -23 -121 23 -109
rect -23 -1097 -17 -121
rect 17 -1097 23 -121
rect -23 -1109 23 -1097
rect 235 -121 281 -109
rect 235 -1097 241 -121
rect 275 -1097 281 -121
rect 235 -1109 281 -1097
rect 493 -121 539 -109
rect 493 -1097 499 -121
rect 533 -1097 539 -121
rect 493 -1109 539 -1097
rect 751 -121 797 -109
rect 751 -1097 757 -121
rect 791 -1097 797 -121
rect 751 -1109 797 -1097
rect 1009 -121 1055 -109
rect 1009 -1097 1015 -121
rect 1049 -1097 1055 -121
rect 1009 -1109 1055 -1097
rect 1267 -121 1313 -109
rect 1267 -1097 1273 -121
rect 1307 -1097 1313 -121
rect 1267 -1109 1313 -1097
rect -1223 -1147 -1099 -1141
rect -1223 -1181 -1211 -1147
rect -1111 -1181 -1099 -1147
rect -1223 -1187 -1099 -1181
rect -965 -1147 -841 -1141
rect -965 -1181 -953 -1147
rect -853 -1181 -841 -1147
rect -965 -1187 -841 -1181
rect -707 -1147 -583 -1141
rect -707 -1181 -695 -1147
rect -595 -1181 -583 -1147
rect -707 -1187 -583 -1181
rect -449 -1147 -325 -1141
rect -449 -1181 -437 -1147
rect -337 -1181 -325 -1147
rect -449 -1187 -325 -1181
rect -191 -1147 -67 -1141
rect -191 -1181 -179 -1147
rect -79 -1181 -67 -1147
rect -191 -1187 -67 -1181
rect 67 -1147 191 -1141
rect 67 -1181 79 -1147
rect 179 -1181 191 -1147
rect 67 -1187 191 -1181
rect 325 -1147 449 -1141
rect 325 -1181 337 -1147
rect 437 -1181 449 -1147
rect 325 -1187 449 -1181
rect 583 -1147 707 -1141
rect 583 -1181 595 -1147
rect 695 -1181 707 -1147
rect 583 -1187 707 -1181
rect 841 -1147 965 -1141
rect 841 -1181 853 -1147
rect 953 -1181 965 -1147
rect 841 -1187 965 -1181
rect 1099 -1147 1223 -1141
rect 1099 -1181 1111 -1147
rect 1211 -1181 1223 -1147
rect 1099 -1187 1223 -1181
<< properties >>
string FIXED_BBOX -1404 -1266 1404 1266
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 5 l 1 m 2 nf 10 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
