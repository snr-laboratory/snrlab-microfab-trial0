magic
tech sky130B
magscale 1 2
timestamp 1686775877
<< nwell >>
rect -2457 -1219 2457 1219
<< pmoslvt >>
rect -2261 -1000 -1861 1000
rect -1803 -1000 -1403 1000
rect -1345 -1000 -945 1000
rect -887 -1000 -487 1000
rect -429 -1000 -29 1000
rect 29 -1000 429 1000
rect 487 -1000 887 1000
rect 945 -1000 1345 1000
rect 1403 -1000 1803 1000
rect 1861 -1000 2261 1000
<< pdiff >>
rect -2319 988 -2261 1000
rect -2319 -988 -2307 988
rect -2273 -988 -2261 988
rect -2319 -1000 -2261 -988
rect -1861 988 -1803 1000
rect -1861 -988 -1849 988
rect -1815 -988 -1803 988
rect -1861 -1000 -1803 -988
rect -1403 988 -1345 1000
rect -1403 -988 -1391 988
rect -1357 -988 -1345 988
rect -1403 -1000 -1345 -988
rect -945 988 -887 1000
rect -945 -988 -933 988
rect -899 -988 -887 988
rect -945 -1000 -887 -988
rect -487 988 -429 1000
rect -487 -988 -475 988
rect -441 -988 -429 988
rect -487 -1000 -429 -988
rect -29 988 29 1000
rect -29 -988 -17 988
rect 17 -988 29 988
rect -29 -1000 29 -988
rect 429 988 487 1000
rect 429 -988 441 988
rect 475 -988 487 988
rect 429 -1000 487 -988
rect 887 988 945 1000
rect 887 -988 899 988
rect 933 -988 945 988
rect 887 -1000 945 -988
rect 1345 988 1403 1000
rect 1345 -988 1357 988
rect 1391 -988 1403 988
rect 1345 -1000 1403 -988
rect 1803 988 1861 1000
rect 1803 -988 1815 988
rect 1849 -988 1861 988
rect 1803 -1000 1861 -988
rect 2261 988 2319 1000
rect 2261 -988 2273 988
rect 2307 -988 2319 988
rect 2261 -1000 2319 -988
<< pdiffc >>
rect -2307 -988 -2273 988
rect -1849 -988 -1815 988
rect -1391 -988 -1357 988
rect -933 -988 -899 988
rect -475 -988 -441 988
rect -17 -988 17 988
rect 441 -988 475 988
rect 899 -988 933 988
rect 1357 -988 1391 988
rect 1815 -988 1849 988
rect 2273 -988 2307 988
<< nsubdiff >>
rect -2421 1149 -2325 1183
rect 2325 1149 2421 1183
rect -2421 1087 -2387 1149
rect 2387 1087 2421 1149
rect -2421 -1149 -2387 -1087
rect 2387 -1149 2421 -1087
rect -2421 -1183 -2325 -1149
rect 2325 -1183 2421 -1149
<< nsubdiffcont >>
rect -2325 1149 2325 1183
rect -2421 -1087 -2387 1087
rect 2387 -1087 2421 1087
rect -2325 -1183 2325 -1149
<< poly >>
rect -2169 1081 -1953 1097
rect -2169 1064 -2153 1081
rect -2261 1047 -2153 1064
rect -1969 1064 -1953 1081
rect -1711 1081 -1495 1097
rect -1711 1064 -1695 1081
rect -1969 1047 -1861 1064
rect -2261 1000 -1861 1047
rect -1803 1047 -1695 1064
rect -1511 1064 -1495 1081
rect -1253 1081 -1037 1097
rect -1253 1064 -1237 1081
rect -1511 1047 -1403 1064
rect -1803 1000 -1403 1047
rect -1345 1047 -1237 1064
rect -1053 1064 -1037 1081
rect -795 1081 -579 1097
rect -795 1064 -779 1081
rect -1053 1047 -945 1064
rect -1345 1000 -945 1047
rect -887 1047 -779 1064
rect -595 1064 -579 1081
rect -337 1081 -121 1097
rect -337 1064 -321 1081
rect -595 1047 -487 1064
rect -887 1000 -487 1047
rect -429 1047 -321 1064
rect -137 1064 -121 1081
rect 121 1081 337 1097
rect 121 1064 137 1081
rect -137 1047 -29 1064
rect -429 1000 -29 1047
rect 29 1047 137 1064
rect 321 1064 337 1081
rect 579 1081 795 1097
rect 579 1064 595 1081
rect 321 1047 429 1064
rect 29 1000 429 1047
rect 487 1047 595 1064
rect 779 1064 795 1081
rect 1037 1081 1253 1097
rect 1037 1064 1053 1081
rect 779 1047 887 1064
rect 487 1000 887 1047
rect 945 1047 1053 1064
rect 1237 1064 1253 1081
rect 1495 1081 1711 1097
rect 1495 1064 1511 1081
rect 1237 1047 1345 1064
rect 945 1000 1345 1047
rect 1403 1047 1511 1064
rect 1695 1064 1711 1081
rect 1953 1081 2169 1097
rect 1953 1064 1969 1081
rect 1695 1047 1803 1064
rect 1403 1000 1803 1047
rect 1861 1047 1969 1064
rect 2153 1064 2169 1081
rect 2153 1047 2261 1064
rect 1861 1000 2261 1047
rect -2261 -1047 -1861 -1000
rect -2261 -1064 -2153 -1047
rect -2169 -1081 -2153 -1064
rect -1969 -1064 -1861 -1047
rect -1803 -1047 -1403 -1000
rect -1803 -1064 -1695 -1047
rect -1969 -1081 -1953 -1064
rect -2169 -1097 -1953 -1081
rect -1711 -1081 -1695 -1064
rect -1511 -1064 -1403 -1047
rect -1345 -1047 -945 -1000
rect -1345 -1064 -1237 -1047
rect -1511 -1081 -1495 -1064
rect -1711 -1097 -1495 -1081
rect -1253 -1081 -1237 -1064
rect -1053 -1064 -945 -1047
rect -887 -1047 -487 -1000
rect -887 -1064 -779 -1047
rect -1053 -1081 -1037 -1064
rect -1253 -1097 -1037 -1081
rect -795 -1081 -779 -1064
rect -595 -1064 -487 -1047
rect -429 -1047 -29 -1000
rect -429 -1064 -321 -1047
rect -595 -1081 -579 -1064
rect -795 -1097 -579 -1081
rect -337 -1081 -321 -1064
rect -137 -1064 -29 -1047
rect 29 -1047 429 -1000
rect 29 -1064 137 -1047
rect -137 -1081 -121 -1064
rect -337 -1097 -121 -1081
rect 121 -1081 137 -1064
rect 321 -1064 429 -1047
rect 487 -1047 887 -1000
rect 487 -1064 595 -1047
rect 321 -1081 337 -1064
rect 121 -1097 337 -1081
rect 579 -1081 595 -1064
rect 779 -1064 887 -1047
rect 945 -1047 1345 -1000
rect 945 -1064 1053 -1047
rect 779 -1081 795 -1064
rect 579 -1097 795 -1081
rect 1037 -1081 1053 -1064
rect 1237 -1064 1345 -1047
rect 1403 -1047 1803 -1000
rect 1403 -1064 1511 -1047
rect 1237 -1081 1253 -1064
rect 1037 -1097 1253 -1081
rect 1495 -1081 1511 -1064
rect 1695 -1064 1803 -1047
rect 1861 -1047 2261 -1000
rect 1861 -1064 1969 -1047
rect 1695 -1081 1711 -1064
rect 1495 -1097 1711 -1081
rect 1953 -1081 1969 -1064
rect 2153 -1064 2261 -1047
rect 2153 -1081 2169 -1064
rect 1953 -1097 2169 -1081
<< polycont >>
rect -2153 1047 -1969 1081
rect -1695 1047 -1511 1081
rect -1237 1047 -1053 1081
rect -779 1047 -595 1081
rect -321 1047 -137 1081
rect 137 1047 321 1081
rect 595 1047 779 1081
rect 1053 1047 1237 1081
rect 1511 1047 1695 1081
rect 1969 1047 2153 1081
rect -2153 -1081 -1969 -1047
rect -1695 -1081 -1511 -1047
rect -1237 -1081 -1053 -1047
rect -779 -1081 -595 -1047
rect -321 -1081 -137 -1047
rect 137 -1081 321 -1047
rect 595 -1081 779 -1047
rect 1053 -1081 1237 -1047
rect 1511 -1081 1695 -1047
rect 1969 -1081 2153 -1047
<< locali >>
rect -2421 1149 -2325 1183
rect 2325 1149 2421 1183
rect -2421 1087 -2387 1149
rect 2387 1087 2421 1149
rect -2169 1047 -2153 1081
rect -1969 1047 -1953 1081
rect -1711 1047 -1695 1081
rect -1511 1047 -1495 1081
rect -1253 1047 -1237 1081
rect -1053 1047 -1037 1081
rect -795 1047 -779 1081
rect -595 1047 -579 1081
rect -337 1047 -321 1081
rect -137 1047 -121 1081
rect 121 1047 137 1081
rect 321 1047 337 1081
rect 579 1047 595 1081
rect 779 1047 795 1081
rect 1037 1047 1053 1081
rect 1237 1047 1253 1081
rect 1495 1047 1511 1081
rect 1695 1047 1711 1081
rect 1953 1047 1969 1081
rect 2153 1047 2169 1081
rect -2307 988 -2273 1004
rect -2307 -1004 -2273 -988
rect -1849 988 -1815 1004
rect -1849 -1004 -1815 -988
rect -1391 988 -1357 1004
rect -1391 -1004 -1357 -988
rect -933 988 -899 1004
rect -933 -1004 -899 -988
rect -475 988 -441 1004
rect -475 -1004 -441 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 441 988 475 1004
rect 441 -1004 475 -988
rect 899 988 933 1004
rect 899 -1004 933 -988
rect 1357 988 1391 1004
rect 1357 -1004 1391 -988
rect 1815 988 1849 1004
rect 1815 -1004 1849 -988
rect 2273 988 2307 1004
rect 2273 -1004 2307 -988
rect -2169 -1081 -2153 -1047
rect -1969 -1081 -1953 -1047
rect -1711 -1081 -1695 -1047
rect -1511 -1081 -1495 -1047
rect -1253 -1081 -1237 -1047
rect -1053 -1081 -1037 -1047
rect -795 -1081 -779 -1047
rect -595 -1081 -579 -1047
rect -337 -1081 -321 -1047
rect -137 -1081 -121 -1047
rect 121 -1081 137 -1047
rect 321 -1081 337 -1047
rect 579 -1081 595 -1047
rect 779 -1081 795 -1047
rect 1037 -1081 1053 -1047
rect 1237 -1081 1253 -1047
rect 1495 -1081 1511 -1047
rect 1695 -1081 1711 -1047
rect 1953 -1081 1969 -1047
rect 2153 -1081 2169 -1047
rect -2421 -1149 -2387 -1087
rect 2387 -1149 2421 -1087
rect -2421 -1183 -2325 -1149
rect 2325 -1183 2421 -1149
<< viali >>
rect -2153 1047 -1969 1081
rect -1695 1047 -1511 1081
rect -1237 1047 -1053 1081
rect -779 1047 -595 1081
rect -321 1047 -137 1081
rect 137 1047 321 1081
rect 595 1047 779 1081
rect 1053 1047 1237 1081
rect 1511 1047 1695 1081
rect 1969 1047 2153 1081
rect -2307 -988 -2273 988
rect -1849 -988 -1815 988
rect -1391 -988 -1357 988
rect -933 -988 -899 988
rect -475 -988 -441 988
rect -17 -988 17 988
rect 441 -988 475 988
rect 899 -988 933 988
rect 1357 -988 1391 988
rect 1815 -988 1849 988
rect 2273 -988 2307 988
rect -2153 -1081 -1969 -1047
rect -1695 -1081 -1511 -1047
rect -1237 -1081 -1053 -1047
rect -779 -1081 -595 -1047
rect -321 -1081 -137 -1047
rect 137 -1081 321 -1047
rect 595 -1081 779 -1047
rect 1053 -1081 1237 -1047
rect 1511 -1081 1695 -1047
rect 1969 -1081 2153 -1047
<< metal1 >>
rect -2165 1081 -1957 1087
rect -2165 1047 -2153 1081
rect -1969 1047 -1957 1081
rect -2165 1041 -1957 1047
rect -1707 1081 -1499 1087
rect -1707 1047 -1695 1081
rect -1511 1047 -1499 1081
rect -1707 1041 -1499 1047
rect -1249 1081 -1041 1087
rect -1249 1047 -1237 1081
rect -1053 1047 -1041 1081
rect -1249 1041 -1041 1047
rect -791 1081 -583 1087
rect -791 1047 -779 1081
rect -595 1047 -583 1081
rect -791 1041 -583 1047
rect -333 1081 -125 1087
rect -333 1047 -321 1081
rect -137 1047 -125 1081
rect -333 1041 -125 1047
rect 125 1081 333 1087
rect 125 1047 137 1081
rect 321 1047 333 1081
rect 125 1041 333 1047
rect 583 1081 791 1087
rect 583 1047 595 1081
rect 779 1047 791 1081
rect 583 1041 791 1047
rect 1041 1081 1249 1087
rect 1041 1047 1053 1081
rect 1237 1047 1249 1081
rect 1041 1041 1249 1047
rect 1499 1081 1707 1087
rect 1499 1047 1511 1081
rect 1695 1047 1707 1081
rect 1499 1041 1707 1047
rect 1957 1081 2165 1087
rect 1957 1047 1969 1081
rect 2153 1047 2165 1081
rect 1957 1041 2165 1047
rect -2313 988 -2267 1000
rect -2313 -988 -2307 988
rect -2273 -988 -2267 988
rect -2313 -1000 -2267 -988
rect -1855 988 -1809 1000
rect -1855 -988 -1849 988
rect -1815 -988 -1809 988
rect -1855 -1000 -1809 -988
rect -1397 988 -1351 1000
rect -1397 -988 -1391 988
rect -1357 -988 -1351 988
rect -1397 -1000 -1351 -988
rect -939 988 -893 1000
rect -939 -988 -933 988
rect -899 -988 -893 988
rect -939 -1000 -893 -988
rect -481 988 -435 1000
rect -481 -988 -475 988
rect -441 -988 -435 988
rect -481 -1000 -435 -988
rect -23 988 23 1000
rect -23 -988 -17 988
rect 17 -988 23 988
rect -23 -1000 23 -988
rect 435 988 481 1000
rect 435 -988 441 988
rect 475 -988 481 988
rect 435 -1000 481 -988
rect 893 988 939 1000
rect 893 -988 899 988
rect 933 -988 939 988
rect 893 -1000 939 -988
rect 1351 988 1397 1000
rect 1351 -988 1357 988
rect 1391 -988 1397 988
rect 1351 -1000 1397 -988
rect 1809 988 1855 1000
rect 1809 -988 1815 988
rect 1849 -988 1855 988
rect 1809 -1000 1855 -988
rect 2267 988 2313 1000
rect 2267 -988 2273 988
rect 2307 -988 2313 988
rect 2267 -1000 2313 -988
rect -2165 -1047 -1957 -1041
rect -2165 -1081 -2153 -1047
rect -1969 -1081 -1957 -1047
rect -2165 -1087 -1957 -1081
rect -1707 -1047 -1499 -1041
rect -1707 -1081 -1695 -1047
rect -1511 -1081 -1499 -1047
rect -1707 -1087 -1499 -1081
rect -1249 -1047 -1041 -1041
rect -1249 -1081 -1237 -1047
rect -1053 -1081 -1041 -1047
rect -1249 -1087 -1041 -1081
rect -791 -1047 -583 -1041
rect -791 -1081 -779 -1047
rect -595 -1081 -583 -1047
rect -791 -1087 -583 -1081
rect -333 -1047 -125 -1041
rect -333 -1081 -321 -1047
rect -137 -1081 -125 -1047
rect -333 -1087 -125 -1081
rect 125 -1047 333 -1041
rect 125 -1081 137 -1047
rect 321 -1081 333 -1047
rect 125 -1087 333 -1081
rect 583 -1047 791 -1041
rect 583 -1081 595 -1047
rect 779 -1081 791 -1047
rect 583 -1087 791 -1081
rect 1041 -1047 1249 -1041
rect 1041 -1081 1053 -1047
rect 1237 -1081 1249 -1047
rect 1041 -1087 1249 -1081
rect 1499 -1047 1707 -1041
rect 1499 -1081 1511 -1047
rect 1695 -1081 1707 -1047
rect 1499 -1087 1707 -1081
rect 1957 -1047 2165 -1041
rect 1957 -1081 1969 -1047
rect 2153 -1081 2165 -1047
rect 1957 -1087 2165 -1081
<< properties >>
string FIXED_BBOX -2404 -1166 2404 1166
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 10 l 2 m 1 nf 10 diffcov 100 polycov 50 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
