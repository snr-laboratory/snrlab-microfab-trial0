magic
tech sky130B
magscale 1 2
timestamp 1686778814
<< nwell >>
rect 1358 2252 1364 2340
<< locali >>
rect -984 5664 8240 5676
rect -984 5364 -972 5664
rect 8226 5364 8240 5664
rect -984 5284 8240 5364
rect -984 2982 -218 5284
rect 422 4490 1704 5284
rect 2206 4490 3400 5284
rect 422 2982 1296 4490
rect -984 2472 1296 2982
rect 2628 2960 3400 4490
rect -298 2466 1296 2472
rect 422 2146 1296 2466
rect 3254 1198 3400 2502
rect 626 150 3400 1198
rect 626 -316 976 150
rect 3254 -316 3400 150
rect 5672 -316 5890 2510
rect -998 -328 8250 -316
rect -998 -864 -986 -328
rect 8238 -864 8250 -328
rect -998 -876 8250 -864
<< viali >>
rect -972 5364 8226 5664
rect -986 -864 8238 -328
<< metal1 >>
rect -984 5664 8240 5676
rect -984 5364 -972 5664
rect 8226 5364 8240 5664
rect -984 5352 8240 5364
rect -292 3132 -104 5352
rect 1858 5208 2056 5352
rect -8 5102 350 5196
rect 1784 5102 3292 5110
rect -8 5100 3292 5102
rect -8 5078 3184 5100
rect -8 4824 12 5078
rect 278 4824 3184 5078
rect -8 4812 3184 4824
rect 3290 4812 3300 5100
rect -8 4802 3292 4812
rect -8 3096 350 4802
rect 1846 4730 2070 4752
rect 1816 4458 2102 4730
rect 1494 4382 1738 4384
rect -36 3066 350 3096
rect 802 2815 1364 4340
rect -690 2593 1364 2815
rect -980 324 -836 2322
rect -690 274 -468 2593
rect -332 -316 -150 2324
rect 6 2290 194 2366
rect 6 1940 14 2290
rect 186 1940 194 2290
rect 6 276 194 1940
rect 354 64 536 2324
rect 802 1704 1364 2593
rect 1472 4330 1756 4382
rect 1842 4354 2074 4458
rect 1472 2388 1526 4330
rect 1708 2388 1756 4330
rect 1472 2292 1756 2388
rect 1816 4352 2074 4354
rect 1816 2578 2102 4352
rect 1816 2356 1846 2578
rect 2074 2356 2102 2578
rect 1816 2340 2102 2356
rect 2160 4332 2444 4394
rect 2160 2390 2214 4332
rect 2396 2390 2444 4332
rect 2160 2332 2444 2390
rect 2152 2296 2444 2332
rect 2554 2296 3116 4340
rect 3426 3134 3562 5352
rect 3608 3094 3618 5174
rect 3826 3094 3836 5174
rect 3608 3092 3836 3094
rect 3880 2914 4016 5134
rect 4066 3094 4076 5174
rect 4284 3094 4294 5174
rect 4338 3134 4474 5352
rect 4066 3092 4294 3094
rect 4524 3094 4534 5174
rect 4742 3094 4752 5174
rect 4524 3092 4752 3094
rect 4800 2914 4936 5134
rect 4982 3094 4992 5174
rect 5200 3094 5210 5174
rect 5256 3132 5392 5352
rect 4982 3092 5210 3094
rect 5440 3094 5450 5174
rect 5658 3094 5668 5174
rect 5440 3092 5668 3094
rect 5714 2914 5850 5170
rect 5898 3094 5908 5174
rect 6116 3094 6126 5174
rect 6174 3132 6310 5352
rect 5898 3092 6126 3094
rect 6356 3094 6366 5174
rect 6574 3094 6584 5174
rect 6356 3092 6584 3094
rect 6632 2914 6768 5170
rect 6814 3094 6824 5174
rect 7032 3094 7042 5174
rect 7088 3132 7224 5352
rect 6814 3092 7042 3094
rect 7272 3094 7282 5174
rect 7490 3094 7500 5174
rect 7272 3092 7500 3094
rect 7548 2914 7684 5170
rect 7730 3094 7740 5174
rect 7948 3094 7958 5174
rect 7730 3092 7958 3094
rect 2554 1930 2804 2296
rect 3064 1930 3116 2296
rect 2554 1704 3116 1930
rect 802 1530 2044 1704
rect 2116 1530 3116 1704
rect 3290 2898 7684 2914
rect 3290 2726 7480 2898
rect 7668 2726 7684 2898
rect 3290 2710 7684 2726
rect 3290 2410 3400 2710
rect 8002 2538 8240 5352
rect 3290 2348 5536 2410
rect 3290 1894 3400 2348
rect 3458 2188 3536 2296
rect 5536 2188 5614 2296
rect 5652 2146 5762 2400
rect 3488 2084 5762 2146
rect 5800 2388 5910 2400
rect 8138 2394 8240 2538
rect 5800 2144 5812 2388
rect 3458 1930 3536 2038
rect 5536 1930 5614 2038
rect 3290 1832 5536 1894
rect 1802 1524 2044 1530
rect 1834 1520 2044 1524
rect 1834 1496 2084 1520
rect 770 1352 3148 1496
rect 3290 1378 3400 1832
rect 3458 1672 3536 1780
rect 5536 1672 5614 1780
rect 5652 1628 5762 2084
rect 5798 2082 5812 2144
rect 5800 1628 5812 2082
rect 3510 1566 5762 1628
rect 5798 1566 5812 1628
rect 3458 1414 3536 1522
rect 5536 1414 5614 1522
rect 1834 1328 2084 1352
rect 3290 1316 5536 1378
rect -60 46 536 64
rect -60 -224 -42 46
rect 518 -224 536 46
rect -60 -242 536 -224
rect 626 1030 3116 1276
rect 626 -316 976 1030
rect 3290 862 3400 1316
rect 3458 1156 3536 1264
rect 5536 1156 5614 1264
rect 5652 1112 5762 1566
rect 5800 1112 5812 1566
rect 3510 1050 5762 1112
rect 5798 1050 5812 1112
rect 3458 898 3536 1006
rect 5536 898 5614 1006
rect 3290 800 5536 862
rect 1124 338 3106 358
rect 1124 84 1140 338
rect 3088 84 3106 338
rect 1124 68 3106 84
rect 3290 346 3400 800
rect 3458 640 3536 748
rect 5536 640 5614 748
rect 5652 596 5762 1050
rect 5800 596 5812 1050
rect 3510 534 5762 596
rect 5798 534 5812 596
rect 3458 382 3536 490
rect 5536 382 5614 490
rect 3290 284 5536 346
rect 1084 -36 3150 -26
rect 1084 -126 1838 -36
rect 2082 -126 3150 -36
rect 1084 -134 3150 -126
rect 3290 -170 3400 284
rect 3458 124 3536 232
rect 5536 124 5614 232
rect 5652 80 5762 534
rect 5800 80 5812 534
rect 3510 18 5762 80
rect 5798 30 5812 80
rect 5898 2144 5910 2388
rect 6030 2348 8240 2394
rect 5898 2082 8050 2144
rect 5898 1628 5910 2082
rect 8138 1878 8240 2348
rect 6030 1832 8240 1878
rect 5898 1566 8050 1628
rect 5898 1112 5910 1566
rect 8138 1362 8240 1832
rect 6030 1316 8240 1362
rect 5898 1050 8050 1112
rect 5898 596 5910 1050
rect 8138 846 8240 1316
rect 6030 800 8240 846
rect 5898 534 8050 596
rect 5898 80 5910 534
rect 8138 330 8240 800
rect 6030 284 8240 330
rect 5898 30 8050 80
rect 5798 18 8050 30
rect 3458 -134 3536 -26
rect 5536 -134 5614 -26
rect 1118 -232 1128 -198
rect 1116 -276 1128 -232
rect 3104 -232 3114 -198
rect 3290 -232 5536 -170
rect 3104 -276 3116 -232
rect 1116 -288 3116 -276
rect 5652 -316 5762 18
rect 5988 -134 5998 -26
rect 8062 -134 8072 -26
rect 8138 -186 8240 284
rect 6030 -232 8240 -186
rect -998 -328 8250 -316
rect -998 -864 -986 -328
rect 8238 -864 8250 -328
rect -998 -876 8250 -864
<< via1 >>
rect 2608 5378 3080 5660
rect 12 4824 278 5078
rect 3184 4812 3290 5100
rect 14 1940 186 2290
rect 1526 2388 1708 4330
rect 1846 2356 2074 2578
rect 2214 2390 2396 4332
rect 3618 3094 3826 5176
rect 4076 3094 4284 5176
rect 4534 3094 4742 5176
rect 4992 3094 5200 5176
rect 5450 3094 5658 5176
rect 5908 3094 6116 5176
rect 6366 3094 6574 5176
rect 6824 3094 7032 5176
rect 7282 3094 7490 5176
rect 7740 3094 7948 5176
rect 2804 1930 3064 2296
rect 7480 2726 7668 2898
rect 3536 2188 5536 2296
rect 3536 1930 5536 2038
rect 3536 1672 5536 1780
rect 3536 1414 5536 1522
rect -42 -224 518 46
rect 3536 1156 5536 1264
rect 3536 898 5536 1006
rect 1140 84 3088 338
rect 3536 640 5536 748
rect 3536 382 5536 490
rect 1838 -126 2082 -36
rect 3536 124 5536 232
rect 5812 30 5898 2388
rect 5998 2188 8062 2296
rect 5998 1930 8062 2038
rect 5998 1672 8062 1780
rect 5998 1414 8062 1522
rect 5998 1156 8062 1264
rect 5998 898 8062 1006
rect 5998 640 8062 748
rect 5998 382 8062 490
rect 5998 124 8062 232
rect 3536 -134 5536 -26
rect 1128 -276 3104 -198
rect 5998 -134 8062 -26
<< metal2 >>
rect 2608 5660 3080 5670
rect 2608 5368 3080 5378
rect 3618 5176 3826 5184
rect -984 5078 302 5102
rect -984 4824 12 5078
rect 278 4824 302 5078
rect -984 4802 302 4824
rect 3176 5100 3618 5110
rect 3176 4812 3184 5100
rect 3290 4812 3618 5100
rect 3176 4802 3618 4812
rect 1526 4330 1708 4340
rect 2214 4332 2396 4342
rect 1526 2378 1708 2388
rect 1846 2578 2074 2588
rect 4076 5176 4284 5184
rect 3826 4802 4076 5110
rect 3618 3082 3826 3094
rect 4534 5176 4742 5184
rect 4284 4802 4534 5110
rect 4076 3082 4284 3094
rect 4992 5176 5200 5184
rect 4742 4802 4992 5110
rect 4534 3082 4742 3094
rect 5450 5176 5658 5184
rect 5200 4802 5450 5110
rect 4992 3082 5200 3094
rect 5908 5176 6116 5184
rect 5658 4802 5908 5110
rect 5450 3082 5658 3094
rect 6366 5176 6574 5184
rect 6116 4802 6366 5110
rect 5908 3082 6116 3094
rect 6824 5176 7032 5184
rect 6574 4802 6824 5110
rect 6366 3082 6574 3094
rect 7282 5176 7490 5184
rect 7032 4802 7282 5110
rect 6824 3082 7032 3094
rect 7740 5176 7948 5184
rect 7490 4802 7740 5110
rect 7282 3082 7490 3094
rect 7740 3082 7948 3094
rect 7464 2898 7684 2914
rect 7464 2726 7480 2898
rect 7668 2726 7684 2898
rect 2214 2380 2396 2390
rect 5812 2388 5898 2398
rect 1846 2346 2074 2356
rect 2804 2298 3064 2306
rect 6 2296 3540 2298
rect 6 2290 2804 2296
rect 6 1940 14 2290
rect 186 1940 2804 2290
rect 6 1930 2804 1940
rect 3064 2188 3536 2296
rect 5536 2188 5614 2296
rect 3064 2038 3540 2188
rect 4354 2038 4708 2188
rect 3064 1930 3536 2038
rect 5536 1930 5614 2038
rect 2804 1920 3064 1930
rect 4354 1780 4708 1930
rect 3458 1672 3536 1780
rect 5536 1672 5614 1780
rect 4354 1522 4708 1672
rect 3458 1414 3536 1522
rect 5536 1414 5614 1522
rect 4354 1264 4708 1414
rect 3458 1156 3536 1264
rect 5536 1156 5614 1264
rect 4354 1006 4708 1156
rect 3458 898 3536 1006
rect 5536 898 5614 1006
rect 4354 748 4708 898
rect 3458 640 3536 748
rect 5536 640 5614 748
rect 4354 490 4708 640
rect 3458 382 3536 490
rect 5536 382 5614 490
rect 1140 338 3088 348
rect 4354 232 4708 382
rect 3458 124 3536 232
rect 5536 124 5614 232
rect 1140 74 3088 84
rect -980 46 518 56
rect -980 -224 -42 46
rect 4354 -16 4708 124
rect 7464 2306 7684 2726
rect 5998 2296 8062 2306
rect 5998 2178 8062 2188
rect 6854 2048 7202 2178
rect 5998 2038 8062 2048
rect 5998 1920 8062 1930
rect 6854 1790 7202 1920
rect 5998 1780 8062 1790
rect 5998 1662 8062 1672
rect 6854 1532 7202 1662
rect 5998 1522 8062 1532
rect 5998 1404 8062 1414
rect 6854 1274 7202 1404
rect 5998 1264 8062 1274
rect 5998 1146 8062 1156
rect 6854 1016 7202 1146
rect 5998 1006 8062 1016
rect 5998 888 8062 898
rect 6854 758 7202 888
rect 5998 748 8062 758
rect 5998 630 8062 640
rect 6854 500 7202 630
rect 5998 490 8062 500
rect 5998 372 8062 382
rect 6854 242 7202 372
rect 5998 232 8062 242
rect 5998 114 8062 124
rect 3536 -26 5536 -16
rect 1838 -36 2082 -26
rect 1838 -136 2082 -126
rect 5536 -134 5614 -26
rect 3536 -144 5536 -134
rect -980 -234 518 -224
rect 1128 -198 3104 -188
rect -980 -236 -42 -234
rect 1128 -286 3104 -276
rect 5812 -876 5898 30
rect 6854 -16 7202 114
rect 5998 -26 8062 -16
rect 5998 -144 8062 -134
<< via2 >>
rect 2608 5378 3080 5660
rect 1846 2356 2074 2578
rect 2610 100 3074 324
rect 1838 -126 2082 -36
<< metal3 >>
rect 2588 5660 3090 5676
rect 2588 5378 2608 5660
rect 3080 5378 3090 5660
rect 1828 2578 2090 2592
rect 1828 2356 1846 2578
rect 2074 2356 2090 2578
rect 1828 -31 2090 2356
rect 2588 324 3090 5378
rect 2588 100 2610 324
rect 3074 100 3090 324
rect 2588 74 3090 100
rect 1828 -36 2092 -31
rect 1828 -126 1838 -36
rect 2082 -126 2092 -36
rect 1828 -131 2092 -126
rect 1828 -136 2090 -131
use sky130_fd_pr__pfet_01v8_lvt_JNDTZ3  XM1
timestamp 1686777254
transform 0 1 1957 -1 0 4957
box -396 -319 396 319
use sky130_fd_pr__pfet_01v8_lvt_RHT9FL  XM2
timestamp 1686777254
transform 1 0 1616 0 1 3342
box -396 -1219 396 1219
use sky130_fd_pr__pfet_01v8_lvt_RHT9FL  XM3
timestamp 1686777254
transform -1 0 2302 0 1 3342
box -396 -1219 396 1219
use sky130_fd_pr__nfet_01v8_lvt_MMMA4V  XM4
timestamp 1686775877
transform 0 1 1302 -1 0 1424
box -296 -710 296 710
use sky130_fd_pr__nfet_01v8_lvt_MMMA4V  XM5
timestamp 1686775877
transform 0 1 2616 -1 0 1424
box -296 -710 296 710
use sky130_fd_pr__pfet_01v8_lvt_RHT9FL  XM6
timestamp 1686777254
transform 1 0 102 0 -1 4133
box -396 -1219 396 1219
use sky130_fd_pr__pfet_01v8_lvt_ET3FZ5  XM7
timestamp 1686775877
transform 1 0 5783 0 1 4135
box -2457 -1219 2457 1219
use sky130_fd_pr__nfet_01v8_lvt_JBULW2  XM8
timestamp 1686777446
transform 0 1 4520 -1 0 1081
box -1457 -1210 1457 1210
use sky130_fd_pr__nfet_01v8_lvt_6WXQK8  XM9
timestamp 1686775877
transform 0 1 2116 -1 0 -80
box -296 -1210 296 1210
use sky130_fd_pr__pfet_01v8_lvt_RHT9FL  XM10
timestamp 1686777254
transform 1 0 -584 0 -1 1318
box -396 -1219 396 1219
use sky130_fd_pr__nfet_01v8_lvt_JBULW2  XM11
timestamp 1686777446
transform 0 1 7030 -1 0 1081
box -1457 -1210 1457 1210
use sky130_fd_pr__pfet_01v8_lvt_RHT9FL  XM12
timestamp 1686777254
transform 1 0 102 0 1 1318
box -396 -1219 396 1219
<< labels >>
flabel metal1 -984 5352 -294 5676 0 FreeSans 1024 0 0 0 Vdd
port 1 nsew
flabel metal2 -984 4802 -294 5102 0 FreeSans 1024 0 0 0 Vbp1
port 6 nsew
flabel metal1 -998 -876 -294 -316 0 FreeSans 1024 0 0 0 Vss
port 2 nsew
flabel metal1 -690 2593 -198 2814 0 FreeSans 1024 0 0 0 Vbn1
flabel metal1 2804 2588 3116 2828 0 FreeSans 1024 0 0 0 Vdo
flabel metal2 7480 2726 7668 2898 0 FreeSans 1024 0 0 0 Vbo
port 3 nsew
flabel metal2 5812 -876 5898 -328 0 FreeSans 1024 0 0 0 Vbos
port 10 nsew
flabel metal1 -980 324 -836 2322 0 FreeSans 1024 0 0 0 Vbn1s
port 8 nsew
flabel metal2 -980 -236 -42 56 0 FreeSans 1024 0 0 0 Vdos
port 9 nsew
flabel metal2 1128 -286 3104 -188 0 FreeSans 1024 0 0 0 Vc1s
port 7 nsew
flabel metal3 1828 364 2090 992 0 FreeSans 1024 0 0 0 Vc1
flabel metal2 1526 2388 1708 4330 0 FreeSans 1024 0 0 0 Vinp
port 4 nsew
flabel metal2 2214 2390 2396 4332 0 FreeSans 1024 0 0 0 Vinn
port 5 nsew
<< end >>
