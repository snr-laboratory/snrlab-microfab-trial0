magic
tech sky130B
magscale 1 2
timestamp 1686777446
<< pwell >>
rect -1457 -1210 1457 1210
<< nmoslvt >>
rect -1261 -1000 -1061 1000
rect -1003 -1000 -803 1000
rect -745 -1000 -545 1000
rect -487 -1000 -287 1000
rect -229 -1000 -29 1000
rect 29 -1000 229 1000
rect 287 -1000 487 1000
rect 545 -1000 745 1000
rect 803 -1000 1003 1000
rect 1061 -1000 1261 1000
<< ndiff >>
rect -1319 988 -1261 1000
rect -1319 -988 -1307 988
rect -1273 -988 -1261 988
rect -1319 -1000 -1261 -988
rect -1061 988 -1003 1000
rect -1061 -988 -1049 988
rect -1015 -988 -1003 988
rect -1061 -1000 -1003 -988
rect -803 988 -745 1000
rect -803 -988 -791 988
rect -757 -988 -745 988
rect -803 -1000 -745 -988
rect -545 988 -487 1000
rect -545 -988 -533 988
rect -499 -988 -487 988
rect -545 -1000 -487 -988
rect -287 988 -229 1000
rect -287 -988 -275 988
rect -241 -988 -229 988
rect -287 -1000 -229 -988
rect -29 988 29 1000
rect -29 -988 -17 988
rect 17 -988 29 988
rect -29 -1000 29 -988
rect 229 988 287 1000
rect 229 -988 241 988
rect 275 -988 287 988
rect 229 -1000 287 -988
rect 487 988 545 1000
rect 487 -988 499 988
rect 533 -988 545 988
rect 487 -1000 545 -988
rect 745 988 803 1000
rect 745 -988 757 988
rect 791 -988 803 988
rect 745 -1000 803 -988
rect 1003 988 1061 1000
rect 1003 -988 1015 988
rect 1049 -988 1061 988
rect 1003 -1000 1061 -988
rect 1261 988 1319 1000
rect 1261 -988 1273 988
rect 1307 -988 1319 988
rect 1261 -1000 1319 -988
<< ndiffc >>
rect -1307 -988 -1273 988
rect -1049 -988 -1015 988
rect -791 -988 -757 988
rect -533 -988 -499 988
rect -275 -988 -241 988
rect -17 -988 17 988
rect 241 -988 275 988
rect 499 -988 533 988
rect 757 -988 791 988
rect 1015 -988 1049 988
rect 1273 -988 1307 988
<< psubdiff >>
rect -1421 1140 -1325 1174
rect 1325 1140 1421 1174
rect -1421 1078 -1387 1140
rect 1387 1078 1421 1140
rect -1421 -1140 -1387 -1078
rect 1387 -1140 1421 -1078
rect -1421 -1174 -1325 -1140
rect 1325 -1174 1421 -1140
<< psubdiffcont >>
rect -1325 1140 1325 1174
rect -1421 -1078 -1387 1078
rect 1387 -1078 1421 1078
rect -1325 -1174 1325 -1140
<< poly >>
rect -1219 1072 -1103 1088
rect -1219 1055 -1203 1072
rect -1261 1038 -1203 1055
rect -1119 1055 -1103 1072
rect -961 1072 -845 1088
rect -961 1055 -945 1072
rect -1119 1038 -1061 1055
rect -1261 1000 -1061 1038
rect -1003 1038 -945 1055
rect -861 1055 -845 1072
rect -703 1072 -587 1088
rect -703 1055 -687 1072
rect -861 1038 -803 1055
rect -1003 1000 -803 1038
rect -745 1038 -687 1055
rect -603 1055 -587 1072
rect -445 1072 -329 1088
rect -445 1055 -429 1072
rect -603 1038 -545 1055
rect -745 1000 -545 1038
rect -487 1038 -429 1055
rect -345 1055 -329 1072
rect -187 1072 -71 1088
rect -187 1055 -171 1072
rect -345 1038 -287 1055
rect -487 1000 -287 1038
rect -229 1038 -171 1055
rect -87 1055 -71 1072
rect 71 1072 187 1088
rect 71 1055 87 1072
rect -87 1038 -29 1055
rect -229 1000 -29 1038
rect 29 1038 87 1055
rect 171 1055 187 1072
rect 329 1072 445 1088
rect 329 1055 345 1072
rect 171 1038 229 1055
rect 29 1000 229 1038
rect 287 1038 345 1055
rect 429 1055 445 1072
rect 587 1072 703 1088
rect 587 1055 603 1072
rect 429 1038 487 1055
rect 287 1000 487 1038
rect 545 1038 603 1055
rect 687 1055 703 1072
rect 845 1072 961 1088
rect 845 1055 861 1072
rect 687 1038 745 1055
rect 545 1000 745 1038
rect 803 1038 861 1055
rect 945 1055 961 1072
rect 1103 1072 1219 1088
rect 1103 1055 1119 1072
rect 945 1038 1003 1055
rect 803 1000 1003 1038
rect 1061 1038 1119 1055
rect 1203 1055 1219 1072
rect 1203 1038 1261 1055
rect 1061 1000 1261 1038
rect -1261 -1038 -1061 -1000
rect -1261 -1055 -1203 -1038
rect -1219 -1072 -1203 -1055
rect -1119 -1055 -1061 -1038
rect -1003 -1038 -803 -1000
rect -1003 -1055 -945 -1038
rect -1119 -1072 -1103 -1055
rect -1219 -1088 -1103 -1072
rect -961 -1072 -945 -1055
rect -861 -1055 -803 -1038
rect -745 -1038 -545 -1000
rect -745 -1055 -687 -1038
rect -861 -1072 -845 -1055
rect -961 -1088 -845 -1072
rect -703 -1072 -687 -1055
rect -603 -1055 -545 -1038
rect -487 -1038 -287 -1000
rect -487 -1055 -429 -1038
rect -603 -1072 -587 -1055
rect -703 -1088 -587 -1072
rect -445 -1072 -429 -1055
rect -345 -1055 -287 -1038
rect -229 -1038 -29 -1000
rect -229 -1055 -171 -1038
rect -345 -1072 -329 -1055
rect -445 -1088 -329 -1072
rect -187 -1072 -171 -1055
rect -87 -1055 -29 -1038
rect 29 -1038 229 -1000
rect 29 -1055 87 -1038
rect -87 -1072 -71 -1055
rect -187 -1088 -71 -1072
rect 71 -1072 87 -1055
rect 171 -1055 229 -1038
rect 287 -1038 487 -1000
rect 287 -1055 345 -1038
rect 171 -1072 187 -1055
rect 71 -1088 187 -1072
rect 329 -1072 345 -1055
rect 429 -1055 487 -1038
rect 545 -1038 745 -1000
rect 545 -1055 603 -1038
rect 429 -1072 445 -1055
rect 329 -1088 445 -1072
rect 587 -1072 603 -1055
rect 687 -1055 745 -1038
rect 803 -1038 1003 -1000
rect 803 -1055 861 -1038
rect 687 -1072 703 -1055
rect 587 -1088 703 -1072
rect 845 -1072 861 -1055
rect 945 -1055 1003 -1038
rect 1061 -1038 1261 -1000
rect 1061 -1055 1119 -1038
rect 945 -1072 961 -1055
rect 845 -1088 961 -1072
rect 1103 -1072 1119 -1055
rect 1203 -1055 1261 -1038
rect 1203 -1072 1219 -1055
rect 1103 -1088 1219 -1072
<< polycont >>
rect -1203 1038 -1119 1072
rect -945 1038 -861 1072
rect -687 1038 -603 1072
rect -429 1038 -345 1072
rect -171 1038 -87 1072
rect 87 1038 171 1072
rect 345 1038 429 1072
rect 603 1038 687 1072
rect 861 1038 945 1072
rect 1119 1038 1203 1072
rect -1203 -1072 -1119 -1038
rect -945 -1072 -861 -1038
rect -687 -1072 -603 -1038
rect -429 -1072 -345 -1038
rect -171 -1072 -87 -1038
rect 87 -1072 171 -1038
rect 345 -1072 429 -1038
rect 603 -1072 687 -1038
rect 861 -1072 945 -1038
rect 1119 -1072 1203 -1038
<< locali >>
rect -1421 1140 -1325 1174
rect 1325 1140 1421 1174
rect -1421 1078 -1387 1140
rect 1387 1078 1421 1140
rect -1219 1038 -1203 1072
rect -1119 1038 -1103 1072
rect -961 1038 -945 1072
rect -861 1038 -845 1072
rect -703 1038 -687 1072
rect -603 1038 -587 1072
rect -445 1038 -429 1072
rect -345 1038 -329 1072
rect -187 1038 -171 1072
rect -87 1038 -71 1072
rect 71 1038 87 1072
rect 171 1038 187 1072
rect 329 1038 345 1072
rect 429 1038 445 1072
rect 587 1038 603 1072
rect 687 1038 703 1072
rect 845 1038 861 1072
rect 945 1038 961 1072
rect 1103 1038 1119 1072
rect 1203 1038 1219 1072
rect -1307 988 -1273 1004
rect -1307 -1004 -1273 -988
rect -1049 988 -1015 1004
rect -1049 -1004 -1015 -988
rect -791 988 -757 1004
rect -791 -1004 -757 -988
rect -533 988 -499 1004
rect -533 -1004 -499 -988
rect -275 988 -241 1004
rect -275 -1004 -241 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 241 988 275 1004
rect 241 -1004 275 -988
rect 499 988 533 1004
rect 499 -1004 533 -988
rect 757 988 791 1004
rect 757 -1004 791 -988
rect 1015 988 1049 1004
rect 1015 -1004 1049 -988
rect 1273 988 1307 1004
rect 1273 -1004 1307 -988
rect -1219 -1072 -1203 -1038
rect -1119 -1072 -1103 -1038
rect -961 -1072 -945 -1038
rect -861 -1072 -845 -1038
rect -703 -1072 -687 -1038
rect -603 -1072 -587 -1038
rect -445 -1072 -429 -1038
rect -345 -1072 -329 -1038
rect -187 -1072 -171 -1038
rect -87 -1072 -71 -1038
rect 71 -1072 87 -1038
rect 171 -1072 187 -1038
rect 329 -1072 345 -1038
rect 429 -1072 445 -1038
rect 587 -1072 603 -1038
rect 687 -1072 703 -1038
rect 845 -1072 861 -1038
rect 945 -1072 961 -1038
rect 1103 -1072 1119 -1038
rect 1203 -1072 1219 -1038
rect -1421 -1140 -1387 -1078
rect 1387 -1140 1421 -1078
rect -1421 -1174 -1325 -1140
rect 1325 -1174 1421 -1140
<< viali >>
rect -1203 1038 -1119 1072
rect -945 1038 -861 1072
rect -687 1038 -603 1072
rect -429 1038 -345 1072
rect -171 1038 -87 1072
rect 87 1038 171 1072
rect 345 1038 429 1072
rect 603 1038 687 1072
rect 861 1038 945 1072
rect 1119 1038 1203 1072
rect -1307 -988 -1273 988
rect -1049 -988 -1015 988
rect -791 -988 -757 988
rect -533 -988 -499 988
rect -275 -988 -241 988
rect -17 -988 17 988
rect 241 -988 275 988
rect 499 -988 533 988
rect 757 -988 791 988
rect 1015 -988 1049 988
rect 1273 -988 1307 988
rect -1203 -1072 -1119 -1038
rect -945 -1072 -861 -1038
rect -687 -1072 -603 -1038
rect -429 -1072 -345 -1038
rect -171 -1072 -87 -1038
rect 87 -1072 171 -1038
rect 345 -1072 429 -1038
rect 603 -1072 687 -1038
rect 861 -1072 945 -1038
rect 1119 -1072 1203 -1038
<< metal1 >>
rect -1215 1072 -1107 1078
rect -1215 1038 -1203 1072
rect -1119 1038 -1107 1072
rect -1215 1032 -1107 1038
rect -957 1072 -849 1078
rect -957 1038 -945 1072
rect -861 1038 -849 1072
rect -957 1032 -849 1038
rect -699 1072 -591 1078
rect -699 1038 -687 1072
rect -603 1038 -591 1072
rect -699 1032 -591 1038
rect -441 1072 -333 1078
rect -441 1038 -429 1072
rect -345 1038 -333 1072
rect -441 1032 -333 1038
rect -183 1072 -75 1078
rect -183 1038 -171 1072
rect -87 1038 -75 1072
rect -183 1032 -75 1038
rect 75 1072 183 1078
rect 75 1038 87 1072
rect 171 1038 183 1072
rect 75 1032 183 1038
rect 333 1072 441 1078
rect 333 1038 345 1072
rect 429 1038 441 1072
rect 333 1032 441 1038
rect 591 1072 699 1078
rect 591 1038 603 1072
rect 687 1038 699 1072
rect 591 1032 699 1038
rect 849 1072 957 1078
rect 849 1038 861 1072
rect 945 1038 957 1072
rect 849 1032 957 1038
rect 1107 1072 1215 1078
rect 1107 1038 1119 1072
rect 1203 1038 1215 1072
rect 1107 1032 1215 1038
rect -1313 988 -1267 1000
rect -1313 -988 -1307 988
rect -1273 -988 -1267 988
rect -1313 -1000 -1267 -988
rect -1055 988 -1009 1000
rect -1055 -988 -1049 988
rect -1015 -988 -1009 988
rect -1055 -1000 -1009 -988
rect -797 988 -751 1000
rect -797 -988 -791 988
rect -757 -988 -751 988
rect -797 -1000 -751 -988
rect -539 988 -493 1000
rect -539 -988 -533 988
rect -499 -988 -493 988
rect -539 -1000 -493 -988
rect -281 988 -235 1000
rect -281 -988 -275 988
rect -241 -988 -235 988
rect -281 -1000 -235 -988
rect -23 988 23 1000
rect -23 -988 -17 988
rect 17 -988 23 988
rect -23 -1000 23 -988
rect 235 988 281 1000
rect 235 -988 241 988
rect 275 -988 281 988
rect 235 -1000 281 -988
rect 493 988 539 1000
rect 493 -988 499 988
rect 533 -988 539 988
rect 493 -1000 539 -988
rect 751 988 797 1000
rect 751 -988 757 988
rect 791 -988 797 988
rect 751 -1000 797 -988
rect 1009 988 1055 1000
rect 1009 -988 1015 988
rect 1049 -988 1055 988
rect 1009 -1000 1055 -988
rect 1267 988 1313 1000
rect 1267 -988 1273 988
rect 1307 -988 1313 988
rect 1267 -1000 1313 -988
rect -1215 -1038 -1107 -1032
rect -1215 -1072 -1203 -1038
rect -1119 -1072 -1107 -1038
rect -1215 -1078 -1107 -1072
rect -957 -1038 -849 -1032
rect -957 -1072 -945 -1038
rect -861 -1072 -849 -1038
rect -957 -1078 -849 -1072
rect -699 -1038 -591 -1032
rect -699 -1072 -687 -1038
rect -603 -1072 -591 -1038
rect -699 -1078 -591 -1072
rect -441 -1038 -333 -1032
rect -441 -1072 -429 -1038
rect -345 -1072 -333 -1038
rect -441 -1078 -333 -1072
rect -183 -1038 -75 -1032
rect -183 -1072 -171 -1038
rect -87 -1072 -75 -1038
rect -183 -1078 -75 -1072
rect 75 -1038 183 -1032
rect 75 -1072 87 -1038
rect 171 -1072 183 -1038
rect 75 -1078 183 -1072
rect 333 -1038 441 -1032
rect 333 -1072 345 -1038
rect 429 -1072 441 -1038
rect 333 -1078 441 -1072
rect 591 -1038 699 -1032
rect 591 -1072 603 -1038
rect 687 -1072 699 -1038
rect 591 -1078 699 -1072
rect 849 -1038 957 -1032
rect 849 -1072 861 -1038
rect 945 -1072 957 -1038
rect 849 -1078 957 -1072
rect 1107 -1038 1215 -1032
rect 1107 -1072 1119 -1038
rect 1203 -1072 1215 -1038
rect 1107 -1078 1215 -1072
<< properties >>
string FIXED_BBOX -1404 -1157 1404 1157
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 10 l 1 m 1 nf 10 diffcov 100 polycov 50 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
