magic
tech sky130B
magscale 1 2
timestamp 1686663767
<< locali >>
rect 548 7470 10036 7496
rect 548 7100 570 7470
rect 10020 7100 10036 7470
rect 548 7052 10036 7100
rect 1950 5732 2022 7052
rect 3520 6046 4306 7052
rect 7004 6274 7920 7052
rect 9286 6274 10036 7052
rect 3520 5732 7004 6046
rect 1950 5660 7004 5732
rect 1950 4674 3000 5660
rect 6986 4698 7160 5218
rect 548 3370 858 4376
rect 4324 4148 7160 4698
rect 2206 4146 7160 4148
rect 2206 3890 5274 4146
rect 4834 3370 5274 3890
rect 6622 3472 7160 4146
rect 6622 3370 10000 3472
rect 548 3350 10000 3370
rect 548 2940 560 3350
rect 10020 2940 10036 3350
rect 548 2926 10036 2940
<< viali >>
rect 570 7100 10020 7470
rect 560 2940 10020 3350
<< metal1 >>
rect 548 7470 10036 7496
rect 548 7100 570 7470
rect 10020 7100 10036 7470
rect 548 7088 10036 7100
rect 550 6940 6820 7088
rect 8108 6948 9460 6970
rect 550 6910 3330 6940
rect 550 4840 620 6910
rect 8108 6900 9334 6948
rect 4406 6834 6870 6850
rect 700 6610 3400 6790
rect 4406 6742 4800 6834
rect 5172 6742 6870 6834
rect 4406 6730 6870 6742
rect 7800 6836 9148 6844
rect 700 6100 770 6610
rect 1770 6360 3400 6610
rect 4510 6450 5470 6650
rect 5840 6450 6800 6650
rect 7800 6490 7808 6836
rect 7876 6742 9148 6836
rect 7876 6584 7882 6742
rect 8094 6634 8104 6692
rect 9104 6634 9114 6692
rect 7876 6490 9148 6584
rect 7800 6482 9148 6490
rect 9322 6430 9334 6900
rect 8110 6376 9334 6430
rect 9444 6900 9460 6948
rect 9444 6376 9462 6900
rect 8110 6360 9462 6376
rect 1770 6240 4420 6360
rect 4440 6240 6870 6360
rect 1770 6100 3400 6240
rect 700 6000 3400 6100
rect 680 5990 3400 6000
rect 4770 6136 5200 6160
rect 4770 6044 4800 6136
rect 5172 6044 5200 6136
rect 680 4940 1850 5990
rect 550 4730 1770 4840
rect 2210 4410 2590 5850
rect 2940 5650 3600 5850
rect 3198 5514 3324 5524
rect 1040 4398 2590 4410
rect 1040 4272 2220 4398
rect 2580 4272 2590 4398
rect 1040 4260 2590 4272
rect 2920 4790 3120 5460
rect 2920 4700 2930 4790
rect 3100 4700 3120 4790
rect 1040 4180 2020 4260
rect 990 4050 2070 4180
rect 1050 3700 1990 3970
rect 2920 3770 3120 4700
rect 3198 4888 3208 5514
rect 3314 4888 3324 5514
rect 3198 4434 3324 4888
rect 3400 3940 3600 5650
rect 3684 5514 3810 5524
rect 3684 4888 3694 5514
rect 3800 4888 3810 5514
rect 3684 4434 3810 4888
rect 3400 3850 3410 3940
rect 3590 3850 3600 3940
rect 3400 3840 3600 3850
rect 3880 4190 4080 5460
rect 4770 5100 5200 6044
rect 6100 5184 6530 6160
rect 9708 6110 9894 7088
rect 7264 6036 9894 6110
rect 6100 5178 7158 5184
rect 6100 5118 7050 5178
rect 7150 5118 7158 5178
rect 6100 5110 7158 5118
rect 6100 5100 6530 5110
rect 4138 4900 6850 5010
rect 4138 4398 4270 4900
rect 4520 4800 5480 4810
rect 4520 4690 4540 4800
rect 5460 4690 5480 4800
rect 4520 4670 5480 4690
rect 6460 4550 6790 4810
rect 4764 4406 6790 4550
rect 4128 4272 4138 4398
rect 4270 4272 4280 4398
rect 4764 4190 4942 4406
rect 3880 4052 4942 4190
rect 3880 3770 4080 4052
rect 5460 4020 6760 4120
rect 5460 4010 6440 4020
rect 5260 3940 6490 3950
rect 5260 3850 5270 3940
rect 5370 3850 6490 3940
rect 5260 3840 6490 3850
rect 990 3560 2070 3700
rect 2100 3560 4700 3700
rect 5260 3670 5340 3840
rect 5480 3800 6420 3810
rect 5480 3720 5490 3800
rect 6410 3720 6420 3800
rect 5480 3710 6420 3720
rect 5260 3560 6490 3670
rect 5460 3510 6430 3530
rect 1040 3370 4650 3480
rect 5460 3430 5480 3510
rect 6410 3500 6440 3510
rect 6620 3500 6760 4020
rect 7264 3650 7314 6036
rect 7386 4786 7454 5900
rect 7386 3608 7454 4720
rect 6410 3430 6760 3500
rect 5460 3410 6760 3430
rect 7520 3480 7570 5860
rect 7644 4786 7712 5900
rect 7644 3608 7712 4720
rect 7780 3650 7830 6036
rect 7902 4786 7970 5900
rect 7902 3608 7970 4720
rect 8036 3480 8086 5860
rect 8160 4786 8228 5900
rect 8160 3608 8228 4720
rect 8296 3650 8346 6036
rect 8418 4786 8486 5900
rect 8418 3608 8486 4720
rect 8552 3480 8602 5860
rect 8676 4786 8744 5900
rect 8676 3608 8744 4720
rect 8812 3650 8862 6036
rect 8934 4786 9002 5900
rect 8934 3608 9002 4720
rect 9068 3480 9118 5860
rect 9192 4786 9260 5900
rect 9192 3608 9260 4720
rect 9328 3650 9378 6036
rect 9450 4786 9518 5900
rect 9450 3608 9518 4720
rect 9584 3480 9634 5860
rect 9708 4786 9776 5900
rect 9708 3608 9776 4720
rect 9844 3650 9894 6036
rect 7520 3412 7532 3480
rect 9626 3412 9636 3480
rect 7520 3400 9634 3412
rect 548 3350 10036 3370
rect 548 2940 560 3350
rect 10020 2940 10036 3350
rect 548 2926 10036 2940
<< via1 >>
rect 5570 7100 6320 7470
rect 4800 6742 5172 6834
rect 770 6100 1770 6610
rect 7808 6490 7876 6836
rect 8104 6634 9104 6692
rect 9334 6376 9444 6948
rect 4800 6044 5172 6136
rect 2220 4272 2580 4398
rect 2930 4700 3100 4790
rect 3208 4888 3314 5514
rect 3694 4888 3800 5514
rect 3410 3850 3590 3940
rect 7050 5118 7150 5178
rect 4540 4690 5460 4800
rect 4138 4272 4270 4398
rect 5270 3850 5370 3940
rect 5490 3720 6410 3800
rect 5480 3430 6410 3510
rect 7386 4720 7454 4786
rect 7644 4720 7712 4786
rect 7902 4720 7970 4786
rect 8160 4720 8228 4786
rect 8418 4720 8486 4786
rect 8676 4720 8744 4786
rect 8934 4720 9002 4786
rect 9192 4720 9260 4786
rect 9450 4720 9518 4786
rect 9708 4720 9776 4786
rect 7532 3412 9626 3480
rect 8382 2942 8790 3350
<< metal2 >>
rect 5550 7470 6340 7500
rect 5550 7100 5570 7470
rect 6320 7100 6340 7470
rect 4770 6834 5202 6850
rect 4770 6742 4800 6834
rect 5172 6742 5202 6834
rect 770 6610 1770 6620
rect 770 6090 1770 6100
rect 4770 6136 5202 6742
rect 4770 6044 4800 6136
rect 5172 6044 5202 6136
rect 4770 6020 5202 6044
rect 3208 5514 3314 5524
rect 3208 4878 3314 4888
rect 3694 5514 3800 5524
rect 3694 4878 3800 4888
rect 4540 4800 5460 4810
rect 2920 4790 4540 4800
rect 2920 4700 2930 4790
rect 3100 4700 4540 4790
rect 2920 4690 4540 4700
rect 4540 4680 5460 4690
rect 2580 4408 4282 4410
rect 2220 4398 4282 4408
rect 2580 4272 4138 4398
rect 4270 4272 4282 4398
rect 2220 4262 4282 4272
rect 2580 4260 4282 4262
rect 3400 3940 5370 3950
rect 3400 3850 3410 3940
rect 3590 3850 5270 3940
rect 3400 3840 5370 3850
rect 5550 3810 6340 7100
rect 9334 6948 9444 6958
rect 7800 6836 7884 6844
rect 7800 6490 7808 6836
rect 7876 6490 7884 6836
rect 8104 6692 9104 6702
rect 8104 6624 9104 6634
rect 7800 6482 7884 6490
rect 9334 6366 9444 6376
rect 7044 5178 7158 5184
rect 7044 5118 7050 5178
rect 7150 5118 7158 5178
rect 7044 4790 7158 5118
rect 7044 4786 9790 4790
rect 7044 4720 7386 4786
rect 7454 4720 7644 4786
rect 7712 4720 7902 4786
rect 7970 4720 8160 4786
rect 8228 4720 8418 4786
rect 8486 4720 8676 4786
rect 8744 4720 8934 4786
rect 9002 4720 9192 4786
rect 9260 4720 9450 4786
rect 9518 4720 9708 4786
rect 9776 4720 9790 4786
rect 7044 4716 9790 4720
rect 5490 3800 6410 3810
rect 5490 3710 6410 3720
rect 5480 3510 6410 3520
rect 5480 3420 6410 3430
rect 7532 3480 9626 3490
rect 7532 3402 9626 3412
rect 8364 3350 8808 3370
rect 8364 2942 8382 3350
rect 8790 2942 8808 3350
rect 8364 2926 8808 2942
<< via2 >>
rect 4546 4690 5452 4796
rect 7810 6492 7874 6834
rect 8104 6634 9104 6692
rect 8382 2942 8790 3350
<< metal3 >>
rect 7746 6844 7882 6846
rect 7746 6834 7884 6844
rect 7746 6492 7810 6834
rect 7874 6492 7884 6834
rect 8094 6692 9114 6697
rect 8094 6634 8104 6692
rect 9104 6634 9114 6692
rect 8094 6629 9114 6634
rect 7746 6482 7884 6492
rect 7746 5738 7882 6482
rect 5456 5734 7882 5738
rect 5212 5568 7882 5734
rect 5212 4810 5456 5568
rect 4540 4796 5460 4810
rect 4540 4690 4546 4796
rect 5452 4690 5460 4796
rect 4540 4680 5460 4690
rect 5212 4678 5456 4680
rect 8364 3350 8808 6629
rect 8364 2942 8382 3350
rect 8790 2942 8808 3350
rect 8364 2926 8808 2942
use sky130_fd_pr__pfet_01v8_lvt_9T37YK  XM1
timestamp 1686588514
transform 0 1 3137 -1 0 6392
box -696 -419 696 419
use sky130_fd_pr__pfet_01v8_lvt_LKL9EP  XM2
timestamp 1686588514
transform 1 0 3260 0 1 4977
box -296 -719 296 719
use sky130_fd_pr__pfet_01v8_lvt_LPWSEP  XM3
timestamp 1686588514
transform 1 0 3746 0 1 4977
box -296 -719 296 719
use sky130_fd_pr__nfet_01v8_lvt_MMMA4V  XM4
timestamp 1686573160
transform 0 1 2846 -1 0 3630
box -296 -710 296 710
use sky130_fd_pr__nfet_01v8_lvt_MMMA4V  XM5
timestamp 1686573160
transform 0 1 4160 -1 0 3630
box -296 -710 296 710
use sky130_fd_pr__nfet_01v8_lvt_MMMA4V  XM6
timestamp 1686573160
transform 0 1 4998 -1 0 4958
box -296 -710 296 710
use sky130_fd_pr__nfet_01v8_lvt_MMMA4V  XM7
timestamp 1686573160
transform 0 1 6312 -1 0 4958
box -296 -710 296 710
use sky130_fd_pr__pfet_01v8_lvt_LKL9EP  XM8
timestamp 1686588514
transform 0 1 4989 -1 0 6306
box -296 -719 296 719
use sky130_fd_pr__pfet_01v8_lvt_LPWSEP  XM9
timestamp 1686588514
transform 0 1 6321 -1 0 6306
box -296 -719 296 719
use sky130_fd_pr__pfet_01v8_lvt_LPWSEP  XM10
timestamp 1686588514
transform 0 1 4989 -1 0 6792
box -296 -719 296 719
use sky130_fd_pr__pfet_01v8_lvt_LKL9EP  XM11
timestamp 1686588514
transform 0 1 6321 -1 0 6792
box -296 -719 296 719
use sky130_fd_pr__pfet_01v8_lvt_HV57YK  XM12
timestamp 1686588514
transform 0 1 2405 -1 0 6392
box -696 -419 696 419
use sky130_fd_pr__nfet_01v8_lvt_MMMA4V  XM13
timestamp 1686573160
transform 0 1 1532 -1 0 4116
box -296 -710 296 710
use sky130_fd_pr__nfet_01v8_lvt_MMMA4V  XM14
timestamp 1686573160
transform 0 1 1532 -1 0 3630
box -296 -710 296 710
use sky130_fd_pr__pfet_01v8_lvt_RNLRNP  XM15
timestamp 1686588514
transform 0 1 1267 -1 0 5863
box -1225 -719 1225 719
use sky130_fd_pr__nfet_01v8_lvt_T2LYQ7  XM16
timestamp 1686588514
transform 1 0 8580 0 1 4754
box -1457 -1319 1457 1319
use sky130_fd_pr__nfet_01v8_lvt_EY4QWC  XM17
timestamp 1686588514
transform 0 1 5948 -1 0 3758
box -425 -710 425 710
use sky130_fd_pr__pfet_01v8_lvt_ZWP3RP  XM18
timestamp 1686588514
transform 0 1 8603 -1 0 6663
box -425 -719 425 719
<< labels >>
flabel metal2 770 6100 1770 6610 0 FreeSans 1920 0 0 0 Vbp1
port 6 nsew
flabel metal2 5480 3430 6410 3510 0 FreeSans 1920 0 0 0 Vc1s
port 7 nsew
flabel metal1 5570 7100 6320 7470 0 FreeSans 1920 0 0 0 Vdd
port 1 nsew
flabel metal2 7532 3412 9626 3480 0 FreeSans 1920 0 0 0 Vdos
port 9 nsew
flabel metal2 7044 4716 7386 4790 0 FreeSans 1920 0 0 0 Vdo
port 3 nsew
flabel metal2 9334 6376 9444 6948 0 FreeSans 1920 0 0 0 Vc2s
port 8 nsew
flabel metal1 8382 2942 8790 3350 0 FreeSans 1920 0 0 0 Vss
port 2 nsew
flabel metal2 3694 4888 3800 5514 0 FreeSans 1440 0 0 0 Vinn
port 5 nsew
flabel metal2 3208 4888 3314 5514 0 FreeSans 1440 0 0 0 Vinp
port 4 nsew
<< end >>
