magic
tech sky130B
magscale 1 2
timestamp 1686588514
<< nwell >>
rect -1225 -719 1225 719
<< pmoslvt >>
rect -1029 -500 -29 500
rect 29 -500 1029 500
<< pdiff >>
rect -1087 488 -1029 500
rect -1087 -488 -1075 488
rect -1041 -488 -1029 488
rect -1087 -500 -1029 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 1029 488 1087 500
rect 1029 -488 1041 488
rect 1075 -488 1087 488
rect 1029 -500 1087 -488
<< pdiffc >>
rect -1075 -488 -1041 488
rect -17 -488 17 488
rect 1041 -488 1075 488
<< nsubdiff >>
rect -1189 649 -1093 683
rect 1093 649 1189 683
rect -1189 587 -1155 649
rect 1155 587 1189 649
rect -1189 -649 -1155 -587
rect 1155 -649 1189 -587
rect -1189 -683 -1093 -649
rect 1093 -683 1189 -649
<< nsubdiffcont >>
rect -1093 649 1093 683
rect -1189 -587 -1155 587
rect 1155 -587 1189 587
rect -1093 -683 1093 -649
<< poly >>
rect -932 581 -126 597
rect -932 564 -916 581
rect -1029 547 -916 564
rect -142 564 -126 581
rect 126 581 932 597
rect 126 564 142 581
rect -142 547 -29 564
rect -1029 500 -29 547
rect 29 547 142 564
rect 916 564 932 581
rect 916 547 1029 564
rect 29 500 1029 547
rect -1029 -547 -29 -500
rect -1029 -564 -916 -547
rect -932 -581 -916 -564
rect -142 -564 -29 -547
rect 29 -547 1029 -500
rect 29 -564 142 -547
rect -142 -581 -126 -564
rect -932 -597 -126 -581
rect 126 -581 142 -564
rect 916 -564 1029 -547
rect 916 -581 932 -564
rect 126 -597 932 -581
<< polycont >>
rect -916 547 -142 581
rect 142 547 916 581
rect -916 -581 -142 -547
rect 142 -581 916 -547
<< locali >>
rect -1189 649 -1093 683
rect 1093 649 1189 683
rect -1189 587 -1155 649
rect 1155 587 1189 649
rect -932 547 -916 581
rect -142 547 -126 581
rect 126 547 142 581
rect 916 547 932 581
rect -1075 488 -1041 504
rect -1075 -504 -1041 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 1041 488 1075 504
rect 1041 -504 1075 -488
rect -932 -581 -916 -547
rect -142 -581 -126 -547
rect 126 -581 142 -547
rect 916 -581 932 -547
rect -1189 -649 -1155 -587
rect 1155 -649 1189 -587
rect -1189 -683 -1093 -649
rect 1093 -683 1189 -649
<< viali >>
rect -916 547 -142 581
rect 142 547 916 581
rect -1075 -488 -1041 488
rect -17 -488 17 488
rect 1041 -488 1075 488
rect -916 -581 -142 -547
rect 142 -581 916 -547
<< metal1 >>
rect -928 581 -130 587
rect -928 547 -916 581
rect -142 547 -130 581
rect -928 541 -130 547
rect 130 581 928 587
rect 130 547 142 581
rect 916 547 928 581
rect 130 541 928 547
rect -1081 488 -1035 500
rect -1081 -488 -1075 488
rect -1041 -488 -1035 488
rect -1081 -500 -1035 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 1035 488 1081 500
rect 1035 -488 1041 488
rect 1075 -488 1081 488
rect 1035 -500 1081 -488
rect -928 -547 -130 -541
rect -928 -581 -916 -547
rect -142 -581 -130 -547
rect -928 -587 -130 -581
rect 130 -547 928 -541
rect 130 -581 142 -547
rect 916 -581 928 -547
rect 130 -587 928 -581
<< properties >>
string FIXED_BBOX -1172 -666 1172 666
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 5 l 5 m 1 nf 2 diffcov 100 polycov 80 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 80 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
